library IEEE;
	use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity or_4 is
  port
    (
        i_A: in  std_logic_vector(03 downto 00);

        o_F: out std_logic
    );
end or_4;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definition --
--------------------------------------------------------------------------------
architecture dataflow of or_4 is
begin

    o_F <= i_A(03) or i_A(02) or i_A(01) or i_A(00);
  
end dataflow;
--------------------------------------------------------------------------------
