library IEEE;
    use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity full_adder is
    port
    (
        i_A         : in std_logic;
        i_B         : in std_logic;
        i_carry_in  : in std_logic;

        o_sum       : out std_logic;
        o_carry_out : out std_logic
    );
end full_adder;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definition --
--------------------------------------------------------------------------------
architecture structure of full_adder is
    --------------------------------------------------------------------------------
	-- Component Definitions --
	--------------------------------------------------------------------------------
    component xorg2 is
        port
        (
            i_A : in std_logic;
            i_B : in std_logic;

            o_F : out std_logic
        );
    end component;

    component andg2 is
        port
        (
            i_A : in std_logic;
            i_B : in std_logic;

            o_F : out std_logic
        );
    end component;
    
    component org2 is
        port
        (
            i_A : in std_logic;
            i_B : in std_logic;

            o_F : out std_logic
        );
    end component;
    --------------------------------------------------------------------------------

    --------------------------------------------------------------------------------
    -- Internal Signal Definitions --
    --------------------------------------------------------------------------------
    signal s_sum_0:   std_logic; -- sum of first half adder
    signal s_carry_0: std_logic; -- carry of first half adder
    signal s_carry_1: std_logic; -- carry of second half adder
    --------------------------------------------------------------------------------

begin
    --------------------------------------------------------------------------------
    -- Logic Level 0 --
    -- Half adder 0
    --------------------------------------------------------------------------------
    XOR_HA_0: xorg2
    port map
    (
        i_A => i_A,
        i_B => i_B,

        o_F => s_sum_0
    );

    AND_HA_0: andg2
    port map
    (
        i_A => i_A,
        i_B => i_B,

        o_F => s_carry_0
    );
    --------------------------------------------------------------------------------


    --------------------------------------------------------------------------------
    -- Logic Level 1 --
    -- Half adder 1
    --------------------------------------------------------------------------------
    XOR_HA_1: xorg2
    port map
    (
        i_A => s_sum_0,
        i_B => i_carry_in,

        o_F => o_sum
    );

    AND_HA_1: andg2
    port map
    (
        i_A => s_sum_0,
        i_B => i_carry_in,

        o_F => s_carry_1
    );
    --------------------------------------------------------------------------------

    --------------------------------------------------------------------------------
    -- Logic Level 2 --
    -- Carry OR
    --------------------------------------------------------------------------------
    
    OR_0: org2
    port map
    (
        i_A => s_carry_0,
        i_B => s_carry_1,

        o_F => o_carry_out
    );
    --------------------------------------------------------------------------------
end structure;
--------------------------------------------------------------------------------