library IEEE;
	use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity and_3 is
  port
    (
        i_A: in  std_logic_vector(02 downto 00);

        o_F: out std_logic
    );
end and_3;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definition --
--------------------------------------------------------------------------------
architecture dataflow of and_3 is
begin

    o_F <= i_A(02) and i_A(01) and i_A(00);
  
end dataflow;
--------------------------------------------------------------------------------
