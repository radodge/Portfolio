library IEEE;
    use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity mux_2t1 is 
    port
    (
        i_S:  in  std_logic;

        i_D0: in  std_logic;
        i_D1: in  std_logic;
  
        o_O:  out std_logic
    );
end mux_2t1;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definitition --
--------------------------------------------------------------------------------
architecture structure of mux_2t1 is
    --------------------------------------------------------------------------------
    -- Component Definitions --
    --------------------------------------------------------------------------------
    component invg is
        port
        (
            i_A: in  std_logic;

            o_F: out std_logic
        );
    end component;

    component andg2 is
        port
        (
            i_A: in  std_logic;
            i_B: in  std_logic;

            o_F: out std_logic
        );
    end component;
    
    component org2 is
        port
        (
            i_A: in  std_logic;
            i_B: in  std_logic;

            o_F: out std_logic
        );
    end component;
    --------------------------------------------------------------------------------


    --------------------------------------------------------------------------------
    -- Internal Signal Definitions --
    --------------------------------------------------------------------------------
    signal s_S_inv: std_logic; -- output of inverter, ~S
    signal s_Y0:    std_logic; -- output of ~S & D0
    signal s_Y1:    std_logic; -- output of S & D1
    --------------------------------------------------------------------------------


begin
    --------------------------------------------------------------------------------
    -- Logic Level 0 --
    --------------------------------------------------------------------------------
    inverter: invg 
        port map
        (
            i_A => i_S,

            o_F => s_S_inv
        );
    --------------------------------------------------------------------------------


    --------------------------------------------------------------------------------
    -- Logic Level 1 --
    --------------------------------------------------------------------------------
    and_0: andg2 
        port map
        (
            i_A => s_S_inv,
            i_B => i_D0,

            o_F => s_Y0
        );

    and_1: andg2 
        port map
        (
            i_A => i_S,
            i_B => i_D1,

            o_F => s_Y1
        );
    --------------------------------------------------------------------------------


    --------------------------------------------------------------------------------
    -- Logic Level 2 --
    --------------------------------------------------------------------------------
    or_0: org2 
        port map
        (
            i_A => s_Y0,
            i_B => s_Y1,

            o_F => o_O
        );
    --------------------------------------------------------------------------------
end structure;
--------------------------------------------------------------------------------