library IEEE;
	use IEEE.std_logic_1164.all;
library work;
    use work.MIPS_types.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity mux_2t1_5 is
	port(
			i_S:  in  std_logic;
			i_D0: in  reg_address;
			i_D1: in  reg_address;
			o_O:  out reg_address
		);
end mux_2t1_5;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definitition --
--------------------------------------------------------------------------------
architecture structural of mux_2t1_5 is
	--------------------------------------------------------------------------------
    -- Component Definitions --
    --------------------------------------------------------------------------------
	component mux_2t1 is
		port
		(
			i_S:  in  std_logic;
			i_D0: in  std_logic;
			i_D1: in  std_logic;
			o_O:  out std_logic
		);
	end component;
	--------------------------------------------------------------------------------
begin
	--------------------------------------------------------------------------------
	-- Generate 32 Instances of mux_2t1 --
	--------------------------------------------------------------------------------
	g_mux_2t1_5: for i in 4 downto 0 
		generate mux_2t1_i: mux_2t1 
			port map
			(
				i_S  => i_S,
				i_D0 => i_D0(i),
				i_D1 => i_D1(i),
				o_O  => o_O(i)
			);
		end generate g_mux_2t1_5;
	--------------------------------------------------------------------------------
end structural;
--------------------------------------------------------------------------------