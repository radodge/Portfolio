library IEEE;
    use IEEE.std_logic_1164.all;
library work;
    use work.MIPS_types.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity ones_comp_32 is
    port
    (
        i_A: in  bus_32;

        o_F: out bus_32
    );  
end ones_comp_32;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definitition --
--------------------------------------------------------------------------------
architecture structure of ones_comp_32 is
    --------------------------------------------------------------------------------
    -- Component Definitions --
    --------------------------------------------------------------------------------
    component invg is
        port
        (
            i_A: in std_logic;

            o_F: out std_logic
        );
    end component;
    --------------------------------------------------------------------------------

begin

        G_invg_i: for i in 31 downto 0 
        generate invg_i: invg 
            port map
            (
                i_A => i_A(i),

                o_F => o_F(i)
            );
        end generate G_invg_i;
end structure;
--------------------------------------------------------------------------------