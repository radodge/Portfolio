library IEEE;
	use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity xnor_2 is
  port
    (
        i_A: in  std_logic;
        i_B: in  std_logic;

        o_F: out std_logic
    );
end xnor_2;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definition --
--------------------------------------------------------------------------------
architecture dataflow of xnor_2 is
begin

    o_F <= not(i_A xor i_B);
  
end dataflow;
--------------------------------------------------------------------------------