library IEEE;
    use IEEE.std_logic_1164.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity inv_N is
    generic
    (
        N: integer := 32
    );
    port
    (
        i_A: in  std_logic_vector(N-1 downto 00);

        o_F: out std_logic_vector(N-1 downto 00)
    );
end inv_N;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definition --
--------------------------------------------------------------------------------
architecture structural of inv_N is
    --------------------------------------------------------------------------------
	-- Component Definitions --
	--------------------------------------------------------------------------------
    component invg is
        port
        (
            i_A: in  std_logic;

            o_F: out std_logic
        );
    end component;
    --------------------------------------------------------------------------------
begin
    --------------------------------------------------------------------------------
    -- Generate N Instances of invg
    --------------------------------------------------------------------------------
    G_NBit_inv: for i in N-1 downto 00
    generate invg_i: invg
        port map
        (
            i_A => i_A(i),

            o_F => o_F(i)
        );
    end generate G_NBit_inv;
end structural;
--------------------------------------------------------------------------------