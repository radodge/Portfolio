library IEEE;
	use IEEE.std_logic_1164.all;
library work;
    use work.MIPS_types.all;

--------------------------------------------------------------------------------
-- Top-level Entity Definition --
--------------------------------------------------------------------------------
entity mux_2t1_32 is
	port(
		i_S:  in  std_logic;
		i_D0: in  bus_32;
		i_D1: in  bus_32;
		o_O:  out bus_32
	);
end mux_2t1_32;
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Architecture Definitition --
--------------------------------------------------------------------------------
architecture structural of mux_2t1_32 is
	--------------------------------------------------------------------------------
    -- Component Definitions --
    --------------------------------------------------------------------------------
	component mux_2t1 is
		port
		(
			i_S:  in  std_logic;
			i_D0: in  std_logic;
			i_D1: in  std_logic;
			o_O:  out std_logic
		);
	end component;
	--------------------------------------------------------------------------------
begin
	--------------------------------------------------------------------------------
	-- Generate 32 Instances of mux_2t1 --
	--------------------------------------------------------------------------------
	G_mux_2t1_32: for i in 31 downto 0 
		generate mux_2t1_i: mux_2t1 
			port map
			(
				i_S  => i_S,
				i_D0 => i_D0(i),
				i_D1 => i_D1(i),
				o_O  => o_O(i)
			);
		end generate G_mux_2t1_32;
	--------------------------------------------------------------------------------
end structural;
--------------------------------------------------------------------------------